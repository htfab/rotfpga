magic
tech sky130A
magscale 1 2
timestamp 1636993897
<< obsli1 >>
rect 1104 2159 176519 177361
<< obsm1 >>
rect 106 2128 177362 177676
<< metal2 >>
rect 754 178863 810 179663
rect 2226 178863 2282 179663
rect 3790 178863 3846 179663
rect 5354 178863 5410 179663
rect 6918 178863 6974 179663
rect 8482 178863 8538 179663
rect 10046 178863 10102 179663
rect 11610 178863 11666 179663
rect 13174 178863 13230 179663
rect 14738 178863 14794 179663
rect 16302 178863 16358 179663
rect 17866 178863 17922 179663
rect 19430 178863 19486 179663
rect 20994 178863 21050 179663
rect 22558 178863 22614 179663
rect 24030 178863 24086 179663
rect 25594 178863 25650 179663
rect 27158 178863 27214 179663
rect 28722 178863 28778 179663
rect 30286 178863 30342 179663
rect 31850 178863 31906 179663
rect 33414 178863 33470 179663
rect 34978 178863 35034 179663
rect 36542 178863 36598 179663
rect 38106 178863 38162 179663
rect 39670 178863 39726 179663
rect 41234 178863 41290 179663
rect 42798 178863 42854 179663
rect 44362 178863 44418 179663
rect 45834 178863 45890 179663
rect 47398 178863 47454 179663
rect 48962 178863 49018 179663
rect 50526 178863 50582 179663
rect 52090 178863 52146 179663
rect 53654 178863 53710 179663
rect 55218 178863 55274 179663
rect 56782 178863 56838 179663
rect 58346 178863 58402 179663
rect 59910 178863 59966 179663
rect 61474 178863 61530 179663
rect 63038 178863 63094 179663
rect 64602 178863 64658 179663
rect 66166 178863 66222 179663
rect 67638 178863 67694 179663
rect 69202 178863 69258 179663
rect 70766 178863 70822 179663
rect 72330 178863 72386 179663
rect 73894 178863 73950 179663
rect 75458 178863 75514 179663
rect 77022 178863 77078 179663
rect 78586 178863 78642 179663
rect 80150 178863 80206 179663
rect 81714 178863 81770 179663
rect 83278 178863 83334 179663
rect 84842 178863 84898 179663
rect 86406 178863 86462 179663
rect 87970 178863 88026 179663
rect 89534 178863 89590 179663
rect 91006 178863 91062 179663
rect 92570 178863 92626 179663
rect 94134 178863 94190 179663
rect 95698 178863 95754 179663
rect 97262 178863 97318 179663
rect 98826 178863 98882 179663
rect 100390 178863 100446 179663
rect 101954 178863 102010 179663
rect 103518 178863 103574 179663
rect 105082 178863 105138 179663
rect 106646 178863 106702 179663
rect 108210 178863 108266 179663
rect 109774 178863 109830 179663
rect 111338 178863 111394 179663
rect 112810 178863 112866 179663
rect 114374 178863 114430 179663
rect 115938 178863 115994 179663
rect 117502 178863 117558 179663
rect 119066 178863 119122 179663
rect 120630 178863 120686 179663
rect 122194 178863 122250 179663
rect 123758 178863 123814 179663
rect 125322 178863 125378 179663
rect 126886 178863 126942 179663
rect 128450 178863 128506 179663
rect 130014 178863 130070 179663
rect 131578 178863 131634 179663
rect 133142 178863 133198 179663
rect 134614 178863 134670 179663
rect 136178 178863 136234 179663
rect 137742 178863 137798 179663
rect 139306 178863 139362 179663
rect 140870 178863 140926 179663
rect 142434 178863 142490 179663
rect 143998 178863 144054 179663
rect 145562 178863 145618 179663
rect 147126 178863 147182 179663
rect 148690 178863 148746 179663
rect 150254 178863 150310 179663
rect 151818 178863 151874 179663
rect 153382 178863 153438 179663
rect 154946 178863 155002 179663
rect 156418 178863 156474 179663
rect 157982 178863 158038 179663
rect 159546 178863 159602 179663
rect 161110 178863 161166 179663
rect 162674 178863 162730 179663
rect 164238 178863 164294 179663
rect 165802 178863 165858 179663
rect 167366 178863 167422 179663
rect 168930 178863 168986 179663
rect 170494 178863 170550 179663
rect 172058 178863 172114 179663
rect 173622 178863 173678 179663
rect 175186 178863 175242 179663
rect 176750 178863 176806 179663
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55494 0 55550 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63774 0 63830 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68098 0 68154 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87234 0 87290 800
rect 87602 0 87658 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102690 0 102746 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123206 0 123262 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135442 0 135498 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152094 0 152150 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156418 0 156474 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160742 0 160798 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 164974 0 165030 800
rect 165342 0 165398 800
rect 165710 0 165766 800
rect 166078 0 166134 800
rect 166446 0 166502 800
rect 166814 0 166870 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 167918 0 167974 800
rect 168286 0 168342 800
rect 168654 0 168710 800
rect 169022 0 169078 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 170034 0 170090 800
rect 170402 0 170458 800
rect 170770 0 170826 800
rect 171138 0 171194 800
rect 171506 0 171562 800
rect 171874 0 171930 800
rect 172242 0 172298 800
rect 172610 0 172666 800
rect 172978 0 173034 800
rect 173346 0 173402 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176198 0 176254 800
rect 176566 0 176622 800
rect 176934 0 176990 800
rect 177302 0 177358 800
<< obsm2 >>
rect 112 178807 698 178863
rect 866 178807 2170 178863
rect 2338 178807 3734 178863
rect 3902 178807 5298 178863
rect 5466 178807 6862 178863
rect 7030 178807 8426 178863
rect 8594 178807 9990 178863
rect 10158 178807 11554 178863
rect 11722 178807 13118 178863
rect 13286 178807 14682 178863
rect 14850 178807 16246 178863
rect 16414 178807 17810 178863
rect 17978 178807 19374 178863
rect 19542 178807 20938 178863
rect 21106 178807 22502 178863
rect 22670 178807 23974 178863
rect 24142 178807 25538 178863
rect 25706 178807 27102 178863
rect 27270 178807 28666 178863
rect 28834 178807 30230 178863
rect 30398 178807 31794 178863
rect 31962 178807 33358 178863
rect 33526 178807 34922 178863
rect 35090 178807 36486 178863
rect 36654 178807 38050 178863
rect 38218 178807 39614 178863
rect 39782 178807 41178 178863
rect 41346 178807 42742 178863
rect 42910 178807 44306 178863
rect 44474 178807 45778 178863
rect 45946 178807 47342 178863
rect 47510 178807 48906 178863
rect 49074 178807 50470 178863
rect 50638 178807 52034 178863
rect 52202 178807 53598 178863
rect 53766 178807 55162 178863
rect 55330 178807 56726 178863
rect 56894 178807 58290 178863
rect 58458 178807 59854 178863
rect 60022 178807 61418 178863
rect 61586 178807 62982 178863
rect 63150 178807 64546 178863
rect 64714 178807 66110 178863
rect 66278 178807 67582 178863
rect 67750 178807 69146 178863
rect 69314 178807 70710 178863
rect 70878 178807 72274 178863
rect 72442 178807 73838 178863
rect 74006 178807 75402 178863
rect 75570 178807 76966 178863
rect 77134 178807 78530 178863
rect 78698 178807 80094 178863
rect 80262 178807 81658 178863
rect 81826 178807 83222 178863
rect 83390 178807 84786 178863
rect 84954 178807 86350 178863
rect 86518 178807 87914 178863
rect 88082 178807 89478 178863
rect 89646 178807 90950 178863
rect 91118 178807 92514 178863
rect 92682 178807 94078 178863
rect 94246 178807 95642 178863
rect 95810 178807 97206 178863
rect 97374 178807 98770 178863
rect 98938 178807 100334 178863
rect 100502 178807 101898 178863
rect 102066 178807 103462 178863
rect 103630 178807 105026 178863
rect 105194 178807 106590 178863
rect 106758 178807 108154 178863
rect 108322 178807 109718 178863
rect 109886 178807 111282 178863
rect 111450 178807 112754 178863
rect 112922 178807 114318 178863
rect 114486 178807 115882 178863
rect 116050 178807 117446 178863
rect 117614 178807 119010 178863
rect 119178 178807 120574 178863
rect 120742 178807 122138 178863
rect 122306 178807 123702 178863
rect 123870 178807 125266 178863
rect 125434 178807 126830 178863
rect 126998 178807 128394 178863
rect 128562 178807 129958 178863
rect 130126 178807 131522 178863
rect 131690 178807 133086 178863
rect 133254 178807 134558 178863
rect 134726 178807 136122 178863
rect 136290 178807 137686 178863
rect 137854 178807 139250 178863
rect 139418 178807 140814 178863
rect 140982 178807 142378 178863
rect 142546 178807 143942 178863
rect 144110 178807 145506 178863
rect 145674 178807 147070 178863
rect 147238 178807 148634 178863
rect 148802 178807 150198 178863
rect 150366 178807 151762 178863
rect 151930 178807 153326 178863
rect 153494 178807 154890 178863
rect 155058 178807 156362 178863
rect 156530 178807 157926 178863
rect 158094 178807 159490 178863
rect 159658 178807 161054 178863
rect 161222 178807 162618 178863
rect 162786 178807 164182 178863
rect 164350 178807 165746 178863
rect 165914 178807 167310 178863
rect 167478 178807 168874 178863
rect 169042 178807 170438 178863
rect 170606 178807 172002 178863
rect 172170 178807 173566 178863
rect 173734 178807 175130 178863
rect 175298 178807 176694 178863
rect 176862 178807 177356 178863
rect 112 856 177356 178807
rect 222 800 330 856
rect 498 800 698 856
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3642 856
rect 3810 800 4010 856
rect 4178 800 4286 856
rect 4454 800 4654 856
rect 4822 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6494 856
rect 6662 800 6862 856
rect 7030 800 7230 856
rect 7398 800 7598 856
rect 7766 800 7966 856
rect 8134 800 8334 856
rect 8502 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9346 856
rect 9514 800 9714 856
rect 9882 800 10082 856
rect 10250 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12658 856
rect 12826 800 12934 856
rect 13102 800 13302 856
rect 13470 800 13670 856
rect 13838 800 14038 856
rect 14206 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16614 856
rect 16782 800 16890 856
rect 17058 800 17258 856
rect 17426 800 17626 856
rect 17794 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18730 856
rect 18898 800 19098 856
rect 19266 800 19466 856
rect 19634 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21214 856
rect 21382 800 21582 856
rect 21750 800 21950 856
rect 22118 800 22318 856
rect 22486 800 22686 856
rect 22854 800 23054 856
rect 23222 800 23422 856
rect 23590 800 23790 856
rect 23958 800 24158 856
rect 24326 800 24526 856
rect 24694 800 24894 856
rect 25062 800 25262 856
rect 25430 800 25538 856
rect 25706 800 25906 856
rect 26074 800 26274 856
rect 26442 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27378 856
rect 27546 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29218 856
rect 29386 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30230 856
rect 30398 800 30598 856
rect 30766 800 30966 856
rect 31134 800 31334 856
rect 31502 800 31702 856
rect 31870 800 32070 856
rect 32238 800 32438 856
rect 32606 800 32806 856
rect 32974 800 33174 856
rect 33342 800 33542 856
rect 33710 800 33818 856
rect 33986 800 34186 856
rect 34354 800 34554 856
rect 34722 800 34922 856
rect 35090 800 35290 856
rect 35458 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39614 856
rect 39782 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41822 856
rect 41990 800 42190 856
rect 42358 800 42466 856
rect 42634 800 42834 856
rect 43002 800 43202 856
rect 43370 800 43570 856
rect 43738 800 43938 856
rect 44106 800 44306 856
rect 44474 800 44674 856
rect 44842 800 45042 856
rect 45210 800 45410 856
rect 45578 800 45778 856
rect 45946 800 46146 856
rect 46314 800 46514 856
rect 46682 800 46790 856
rect 46958 800 47158 856
rect 47326 800 47526 856
rect 47694 800 47894 856
rect 48062 800 48262 856
rect 48430 800 48630 856
rect 48798 800 48998 856
rect 49166 800 49366 856
rect 49534 800 49734 856
rect 49902 800 50102 856
rect 50270 800 50470 856
rect 50638 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51482 856
rect 51650 800 51850 856
rect 52018 800 52218 856
rect 52386 800 52586 856
rect 52754 800 52954 856
rect 53122 800 53322 856
rect 53490 800 53690 856
rect 53858 800 54058 856
rect 54226 800 54426 856
rect 54594 800 54794 856
rect 54962 800 55070 856
rect 55238 800 55438 856
rect 55606 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56542 856
rect 56710 800 56910 856
rect 57078 800 57278 856
rect 57446 800 57646 856
rect 57814 800 58014 856
rect 58182 800 58382 856
rect 58550 800 58750 856
rect 58918 800 59118 856
rect 59286 800 59394 856
rect 59562 800 59762 856
rect 59930 800 60130 856
rect 60298 800 60498 856
rect 60666 800 60866 856
rect 61034 800 61234 856
rect 61402 800 61602 856
rect 61770 800 61970 856
rect 62138 800 62338 856
rect 62506 800 62706 856
rect 62874 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63718 856
rect 63886 800 64086 856
rect 64254 800 64454 856
rect 64622 800 64822 856
rect 64990 800 65190 856
rect 65358 800 65558 856
rect 65726 800 65926 856
rect 66094 800 66294 856
rect 66462 800 66662 856
rect 66830 800 67030 856
rect 67198 800 67398 856
rect 67566 800 67674 856
rect 67842 800 68042 856
rect 68210 800 68410 856
rect 68578 800 68778 856
rect 68946 800 69146 856
rect 69314 800 69514 856
rect 69682 800 69882 856
rect 70050 800 70250 856
rect 70418 800 70618 856
rect 70786 800 70986 856
rect 71154 800 71354 856
rect 71522 800 71722 856
rect 71890 800 71998 856
rect 72166 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73102 856
rect 73270 800 73470 856
rect 73638 800 73838 856
rect 74006 800 74206 856
rect 74374 800 74574 856
rect 74742 800 74942 856
rect 75110 800 75310 856
rect 75478 800 75678 856
rect 75846 800 76046 856
rect 76214 800 76322 856
rect 76490 800 76690 856
rect 76858 800 77058 856
rect 77226 800 77426 856
rect 77594 800 77794 856
rect 77962 800 78162 856
rect 78330 800 78530 856
rect 78698 800 78898 856
rect 79066 800 79266 856
rect 79434 800 79634 856
rect 79802 800 80002 856
rect 80170 800 80370 856
rect 80538 800 80646 856
rect 80814 800 81014 856
rect 81182 800 81382 856
rect 81550 800 81750 856
rect 81918 800 82118 856
rect 82286 800 82486 856
rect 82654 800 82854 856
rect 83022 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83958 856
rect 84126 800 84326 856
rect 84494 800 84602 856
rect 84770 800 84970 856
rect 85138 800 85338 856
rect 85506 800 85706 856
rect 85874 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87178 856
rect 87346 800 87546 856
rect 87714 800 87914 856
rect 88082 800 88282 856
rect 88450 800 88650 856
rect 88818 800 88926 856
rect 89094 800 89294 856
rect 89462 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90398 856
rect 90566 800 90766 856
rect 90934 800 91134 856
rect 91302 800 91502 856
rect 91670 800 91870 856
rect 92038 800 92238 856
rect 92406 800 92606 856
rect 92774 800 92974 856
rect 93142 800 93250 856
rect 93418 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94722 856
rect 94890 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95826 856
rect 95994 800 96194 856
rect 96362 800 96562 856
rect 96730 800 96930 856
rect 97098 800 97206 856
rect 97374 800 97574 856
rect 97742 800 97942 856
rect 98110 800 98310 856
rect 98478 800 98678 856
rect 98846 800 99046 856
rect 99214 800 99414 856
rect 99582 800 99782 856
rect 99950 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101254 856
rect 101422 800 101530 856
rect 101698 800 101898 856
rect 102066 800 102266 856
rect 102434 800 102634 856
rect 102802 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104474 856
rect 104642 800 104842 856
rect 105010 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105854 856
rect 106022 800 106222 856
rect 106390 800 106590 856
rect 106758 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107694 856
rect 107862 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108798 856
rect 108966 800 109166 856
rect 109334 800 109534 856
rect 109702 800 109902 856
rect 110070 800 110178 856
rect 110346 800 110546 856
rect 110714 800 110914 856
rect 111082 800 111282 856
rect 111450 800 111650 856
rect 111818 800 112018 856
rect 112186 800 112386 856
rect 112554 800 112754 856
rect 112922 800 113122 856
rect 113290 800 113490 856
rect 113658 800 113858 856
rect 114026 800 114134 856
rect 114302 800 114502 856
rect 114670 800 114870 856
rect 115038 800 115238 856
rect 115406 800 115606 856
rect 115774 800 115974 856
rect 116142 800 116342 856
rect 116510 800 116710 856
rect 116878 800 117078 856
rect 117246 800 117446 856
rect 117614 800 117814 856
rect 117982 800 118182 856
rect 118350 800 118458 856
rect 118626 800 118826 856
rect 118994 800 119194 856
rect 119362 800 119562 856
rect 119730 800 119930 856
rect 120098 800 120298 856
rect 120466 800 120666 856
rect 120834 800 121034 856
rect 121202 800 121402 856
rect 121570 800 121770 856
rect 121938 800 122138 856
rect 122306 800 122506 856
rect 122674 800 122782 856
rect 122950 800 123150 856
rect 123318 800 123518 856
rect 123686 800 123886 856
rect 124054 800 124254 856
rect 124422 800 124622 856
rect 124790 800 124990 856
rect 125158 800 125358 856
rect 125526 800 125726 856
rect 125894 800 126094 856
rect 126262 800 126462 856
rect 126630 800 126830 856
rect 126998 800 127106 856
rect 127274 800 127474 856
rect 127642 800 127842 856
rect 128010 800 128210 856
rect 128378 800 128578 856
rect 128746 800 128946 856
rect 129114 800 129314 856
rect 129482 800 129682 856
rect 129850 800 130050 856
rect 130218 800 130418 856
rect 130586 800 130786 856
rect 130954 800 131062 856
rect 131230 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132166 856
rect 132334 800 132534 856
rect 132702 800 132902 856
rect 133070 800 133270 856
rect 133438 800 133638 856
rect 133806 800 134006 856
rect 134174 800 134374 856
rect 134542 800 134742 856
rect 134910 800 135110 856
rect 135278 800 135386 856
rect 135554 800 135754 856
rect 135922 800 136122 856
rect 136290 800 136490 856
rect 136658 800 136858 856
rect 137026 800 137226 856
rect 137394 800 137594 856
rect 137762 800 137962 856
rect 138130 800 138330 856
rect 138498 800 138698 856
rect 138866 800 139066 856
rect 139234 800 139434 856
rect 139602 800 139710 856
rect 139878 800 140078 856
rect 140246 800 140446 856
rect 140614 800 140814 856
rect 140982 800 141182 856
rect 141350 800 141550 856
rect 141718 800 141918 856
rect 142086 800 142286 856
rect 142454 800 142654 856
rect 142822 800 143022 856
rect 143190 800 143390 856
rect 143558 800 143758 856
rect 143926 800 144034 856
rect 144202 800 144402 856
rect 144570 800 144770 856
rect 144938 800 145138 856
rect 145306 800 145506 856
rect 145674 800 145874 856
rect 146042 800 146242 856
rect 146410 800 146610 856
rect 146778 800 146978 856
rect 147146 800 147346 856
rect 147514 800 147714 856
rect 147882 800 147990 856
rect 148158 800 148358 856
rect 148526 800 148726 856
rect 148894 800 149094 856
rect 149262 800 149462 856
rect 149630 800 149830 856
rect 149998 800 150198 856
rect 150366 800 150566 856
rect 150734 800 150934 856
rect 151102 800 151302 856
rect 151470 800 151670 856
rect 151838 800 152038 856
rect 152206 800 152314 856
rect 152482 800 152682 856
rect 152850 800 153050 856
rect 153218 800 153418 856
rect 153586 800 153786 856
rect 153954 800 154154 856
rect 154322 800 154522 856
rect 154690 800 154890 856
rect 155058 800 155258 856
rect 155426 800 155626 856
rect 155794 800 155994 856
rect 156162 800 156362 856
rect 156530 800 156638 856
rect 156806 800 157006 856
rect 157174 800 157374 856
rect 157542 800 157742 856
rect 157910 800 158110 856
rect 158278 800 158478 856
rect 158646 800 158846 856
rect 159014 800 159214 856
rect 159382 800 159582 856
rect 159750 800 159950 856
rect 160118 800 160318 856
rect 160486 800 160686 856
rect 160854 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162066 856
rect 162234 800 162434 856
rect 162602 800 162802 856
rect 162970 800 163170 856
rect 163338 800 163538 856
rect 163706 800 163906 856
rect 164074 800 164274 856
rect 164442 800 164642 856
rect 164810 800 164918 856
rect 165086 800 165286 856
rect 165454 800 165654 856
rect 165822 800 166022 856
rect 166190 800 166390 856
rect 166558 800 166758 856
rect 166926 800 167126 856
rect 167294 800 167494 856
rect 167662 800 167862 856
rect 168030 800 168230 856
rect 168398 800 168598 856
rect 168766 800 168966 856
rect 169134 800 169242 856
rect 169410 800 169610 856
rect 169778 800 169978 856
rect 170146 800 170346 856
rect 170514 800 170714 856
rect 170882 800 171082 856
rect 171250 800 171450 856
rect 171618 800 171818 856
rect 171986 800 172186 856
rect 172354 800 172554 856
rect 172722 800 172922 856
rect 173090 800 173290 856
rect 173458 800 173566 856
rect 173734 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175038 856
rect 175206 800 175406 856
rect 175574 800 175774 856
rect 175942 800 176142 856
rect 176310 800 176510 856
rect 176678 800 176878 856
rect 177046 800 177246 856
<< obsm3 >>
rect 4208 2143 173488 177377
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< labels >>
rlabel metal2 s 754 178863 810 179663 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 47398 178863 47454 179663 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 52090 178863 52146 179663 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 56782 178863 56838 179663 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 61474 178863 61530 179663 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 66166 178863 66222 179663 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 70766 178863 70822 179663 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 75458 178863 75514 179663 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 80150 178863 80206 179663 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 84842 178863 84898 179663 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 89534 178863 89590 179663 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5354 178863 5410 179663 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 94134 178863 94190 179663 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 98826 178863 98882 179663 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 103518 178863 103574 179663 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 108210 178863 108266 179663 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 112810 178863 112866 179663 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 117502 178863 117558 179663 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 122194 178863 122250 179663 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 126886 178863 126942 179663 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 131578 178863 131634 179663 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 136178 178863 136234 179663 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10046 178863 10102 179663 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 140870 178863 140926 179663 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 145562 178863 145618 179663 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 150254 178863 150310 179663 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 154946 178863 155002 179663 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 159546 178863 159602 179663 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 164238 178863 164294 179663 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 168930 178863 168986 179663 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 173622 178863 173678 179663 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14738 178863 14794 179663 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19430 178863 19486 179663 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24030 178863 24086 179663 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 28722 178863 28778 179663 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33414 178863 33470 179663 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38106 178863 38162 179663 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 42798 178863 42854 179663 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2226 178863 2282 179663 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 48962 178863 49018 179663 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 53654 178863 53710 179663 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 58346 178863 58402 179663 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 63038 178863 63094 179663 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 67638 178863 67694 179663 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 72330 178863 72386 179663 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 77022 178863 77078 179663 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 81714 178863 81770 179663 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 86406 178863 86462 179663 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 91006 178863 91062 179663 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6918 178863 6974 179663 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 95698 178863 95754 179663 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 100390 178863 100446 179663 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 105082 178863 105138 179663 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 109774 178863 109830 179663 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 114374 178863 114430 179663 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 119066 178863 119122 179663 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 123758 178863 123814 179663 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 128450 178863 128506 179663 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 133142 178863 133198 179663 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 137742 178863 137798 179663 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11610 178863 11666 179663 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 142434 178863 142490 179663 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 147126 178863 147182 179663 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 151818 178863 151874 179663 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 156418 178863 156474 179663 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 161110 178863 161166 179663 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 165802 178863 165858 179663 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 170494 178863 170550 179663 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 175186 178863 175242 179663 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16302 178863 16358 179663 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 20994 178863 21050 179663 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 25594 178863 25650 179663 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30286 178863 30342 179663 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 34978 178863 35034 179663 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 39670 178863 39726 179663 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 44362 178863 44418 179663 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3790 178863 3846 179663 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 50526 178863 50582 179663 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 55218 178863 55274 179663 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 59910 178863 59966 179663 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 64602 178863 64658 179663 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 69202 178863 69258 179663 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 73894 178863 73950 179663 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 78586 178863 78642 179663 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 83278 178863 83334 179663 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 87970 178863 88026 179663 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 92570 178863 92626 179663 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8482 178863 8538 179663 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 97262 178863 97318 179663 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 101954 178863 102010 179663 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 106646 178863 106702 179663 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 111338 178863 111394 179663 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 115938 178863 115994 179663 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 120630 178863 120686 179663 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 125322 178863 125378 179663 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 130014 178863 130070 179663 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 134614 178863 134670 179663 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 139306 178863 139362 179663 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13174 178863 13230 179663 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 143998 178863 144054 179663 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 148690 178863 148746 179663 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 153382 178863 153438 179663 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 157982 178863 158038 179663 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 162674 178863 162730 179663 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 167366 178863 167422 179663 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 172058 178863 172114 179663 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 176750 178863 176806 179663 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 17866 178863 17922 179663 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22558 178863 22614 179663 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27158 178863 27214 179663 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 31850 178863 31906 179663 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 36542 178863 36598 179663 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41234 178863 41290 179663 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 45834 178863 45890 179663 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 150990 0 151046 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 152094 0 152150 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 158534 0 158590 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 160742 0 160798 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 168286 0 168342 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 177519 179663
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 51302200
string GDS_START 281178
<< end >>

