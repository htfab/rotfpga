magic
tech sky130A
magscale 1 2
timestamp 1636992219
<< obsli1 >>
rect 1104 2159 89671 90321
<< obsm1 >>
rect 106 2128 90606 90568
<< metal2 >>
rect 386 92026 442 92826
rect 1122 92026 1178 92826
rect 1950 92026 2006 92826
rect 2686 92026 2742 92826
rect 3514 92026 3570 92826
rect 4342 92026 4398 92826
rect 5078 92026 5134 92826
rect 5906 92026 5962 92826
rect 6734 92026 6790 92826
rect 7470 92026 7526 92826
rect 8298 92026 8354 92826
rect 9126 92026 9182 92826
rect 9862 92026 9918 92826
rect 10690 92026 10746 92826
rect 11518 92026 11574 92826
rect 12254 92026 12310 92826
rect 13082 92026 13138 92826
rect 13910 92026 13966 92826
rect 14646 92026 14702 92826
rect 15474 92026 15530 92826
rect 16210 92026 16266 92826
rect 17038 92026 17094 92826
rect 17866 92026 17922 92826
rect 18602 92026 18658 92826
rect 19430 92026 19486 92826
rect 20258 92026 20314 92826
rect 20994 92026 21050 92826
rect 21822 92026 21878 92826
rect 22650 92026 22706 92826
rect 23386 92026 23442 92826
rect 24214 92026 24270 92826
rect 25042 92026 25098 92826
rect 25778 92026 25834 92826
rect 26606 92026 26662 92826
rect 27434 92026 27490 92826
rect 28170 92026 28226 92826
rect 28998 92026 29054 92826
rect 29826 92026 29882 92826
rect 30562 92026 30618 92826
rect 31390 92026 31446 92826
rect 32126 92026 32182 92826
rect 32954 92026 33010 92826
rect 33782 92026 33838 92826
rect 34518 92026 34574 92826
rect 35346 92026 35402 92826
rect 36174 92026 36230 92826
rect 36910 92026 36966 92826
rect 37738 92026 37794 92826
rect 38566 92026 38622 92826
rect 39302 92026 39358 92826
rect 40130 92026 40186 92826
rect 40958 92026 41014 92826
rect 41694 92026 41750 92826
rect 42522 92026 42578 92826
rect 43350 92026 43406 92826
rect 44086 92026 44142 92826
rect 44914 92026 44970 92826
rect 45742 92026 45798 92826
rect 46478 92026 46534 92826
rect 47306 92026 47362 92826
rect 48042 92026 48098 92826
rect 48870 92026 48926 92826
rect 49698 92026 49754 92826
rect 50434 92026 50490 92826
rect 51262 92026 51318 92826
rect 52090 92026 52146 92826
rect 52826 92026 52882 92826
rect 53654 92026 53710 92826
rect 54482 92026 54538 92826
rect 55218 92026 55274 92826
rect 56046 92026 56102 92826
rect 56874 92026 56930 92826
rect 57610 92026 57666 92826
rect 58438 92026 58494 92826
rect 59266 92026 59322 92826
rect 60002 92026 60058 92826
rect 60830 92026 60886 92826
rect 61566 92026 61622 92826
rect 62394 92026 62450 92826
rect 63222 92026 63278 92826
rect 63958 92026 64014 92826
rect 64786 92026 64842 92826
rect 65614 92026 65670 92826
rect 66350 92026 66406 92826
rect 67178 92026 67234 92826
rect 68006 92026 68062 92826
rect 68742 92026 68798 92826
rect 69570 92026 69626 92826
rect 70398 92026 70454 92826
rect 71134 92026 71190 92826
rect 71962 92026 72018 92826
rect 72790 92026 72846 92826
rect 73526 92026 73582 92826
rect 74354 92026 74410 92826
rect 75182 92026 75238 92826
rect 75918 92026 75974 92826
rect 76746 92026 76802 92826
rect 77482 92026 77538 92826
rect 78310 92026 78366 92826
rect 79138 92026 79194 92826
rect 79874 92026 79930 92826
rect 80702 92026 80758 92826
rect 81530 92026 81586 92826
rect 82266 92026 82322 92826
rect 83094 92026 83150 92826
rect 83922 92026 83978 92826
rect 84658 92026 84714 92826
rect 85486 92026 85542 92826
rect 86314 92026 86370 92826
rect 87050 92026 87106 92826
rect 87878 92026 87934 92826
rect 88706 92026 88762 92826
rect 89442 92026 89498 92826
rect 90270 92026 90326 92826
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3790 0 3846 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7286 0 7342 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90638 0 90694 800
<< obsm2 >>
rect 112 91970 330 92026
rect 498 91970 1066 92026
rect 1234 91970 1894 92026
rect 2062 91970 2630 92026
rect 2798 91970 3458 92026
rect 3626 91970 4286 92026
rect 4454 91970 5022 92026
rect 5190 91970 5850 92026
rect 6018 91970 6678 92026
rect 6846 91970 7414 92026
rect 7582 91970 8242 92026
rect 8410 91970 9070 92026
rect 9238 91970 9806 92026
rect 9974 91970 10634 92026
rect 10802 91970 11462 92026
rect 11630 91970 12198 92026
rect 12366 91970 13026 92026
rect 13194 91970 13854 92026
rect 14022 91970 14590 92026
rect 14758 91970 15418 92026
rect 15586 91970 16154 92026
rect 16322 91970 16982 92026
rect 17150 91970 17810 92026
rect 17978 91970 18546 92026
rect 18714 91970 19374 92026
rect 19542 91970 20202 92026
rect 20370 91970 20938 92026
rect 21106 91970 21766 92026
rect 21934 91970 22594 92026
rect 22762 91970 23330 92026
rect 23498 91970 24158 92026
rect 24326 91970 24986 92026
rect 25154 91970 25722 92026
rect 25890 91970 26550 92026
rect 26718 91970 27378 92026
rect 27546 91970 28114 92026
rect 28282 91970 28942 92026
rect 29110 91970 29770 92026
rect 29938 91970 30506 92026
rect 30674 91970 31334 92026
rect 31502 91970 32070 92026
rect 32238 91970 32898 92026
rect 33066 91970 33726 92026
rect 33894 91970 34462 92026
rect 34630 91970 35290 92026
rect 35458 91970 36118 92026
rect 36286 91970 36854 92026
rect 37022 91970 37682 92026
rect 37850 91970 38510 92026
rect 38678 91970 39246 92026
rect 39414 91970 40074 92026
rect 40242 91970 40902 92026
rect 41070 91970 41638 92026
rect 41806 91970 42466 92026
rect 42634 91970 43294 92026
rect 43462 91970 44030 92026
rect 44198 91970 44858 92026
rect 45026 91970 45686 92026
rect 45854 91970 46422 92026
rect 46590 91970 47250 92026
rect 47418 91970 47986 92026
rect 48154 91970 48814 92026
rect 48982 91970 49642 92026
rect 49810 91970 50378 92026
rect 50546 91970 51206 92026
rect 51374 91970 52034 92026
rect 52202 91970 52770 92026
rect 52938 91970 53598 92026
rect 53766 91970 54426 92026
rect 54594 91970 55162 92026
rect 55330 91970 55990 92026
rect 56158 91970 56818 92026
rect 56986 91970 57554 92026
rect 57722 91970 58382 92026
rect 58550 91970 59210 92026
rect 59378 91970 59946 92026
rect 60114 91970 60774 92026
rect 60942 91970 61510 92026
rect 61678 91970 62338 92026
rect 62506 91970 63166 92026
rect 63334 91970 63902 92026
rect 64070 91970 64730 92026
rect 64898 91970 65558 92026
rect 65726 91970 66294 92026
rect 66462 91970 67122 92026
rect 67290 91970 67950 92026
rect 68118 91970 68686 92026
rect 68854 91970 69514 92026
rect 69682 91970 70342 92026
rect 70510 91970 71078 92026
rect 71246 91970 71906 92026
rect 72074 91970 72734 92026
rect 72902 91970 73470 92026
rect 73638 91970 74298 92026
rect 74466 91970 75126 92026
rect 75294 91970 75862 92026
rect 76030 91970 76690 92026
rect 76858 91970 77426 92026
rect 77594 91970 78254 92026
rect 78422 91970 79082 92026
rect 79250 91970 79818 92026
rect 79986 91970 80646 92026
rect 80814 91970 81474 92026
rect 81642 91970 82210 92026
rect 82378 91970 83038 92026
rect 83206 91970 83866 92026
rect 84034 91970 84602 92026
rect 84770 91970 85430 92026
rect 85598 91970 86258 92026
rect 86426 91970 86994 92026
rect 87162 91970 87822 92026
rect 87990 91970 88650 92026
rect 88818 91970 89386 92026
rect 89554 91970 90214 92026
rect 90382 91970 90680 92026
rect 112 856 90680 91970
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 974 856
rect 1142 800 1158 856
rect 1326 800 1342 856
rect 1510 800 1526 856
rect 1694 800 1710 856
rect 1878 800 1894 856
rect 2062 800 2078 856
rect 2246 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 2998 856
rect 3166 800 3182 856
rect 3350 800 3366 856
rect 3534 800 3550 856
rect 3718 800 3734 856
rect 3902 800 3918 856
rect 4086 800 4102 856
rect 4270 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4838 856
rect 5006 800 5022 856
rect 5190 800 5206 856
rect 5374 800 5390 856
rect 5558 800 5574 856
rect 5742 800 5758 856
rect 5926 800 5942 856
rect 6110 800 6126 856
rect 6294 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7046 856
rect 7214 800 7230 856
rect 7398 800 7414 856
rect 7582 800 7598 856
rect 7766 800 7782 856
rect 7950 800 7966 856
rect 8134 800 8150 856
rect 8318 800 8334 856
rect 8502 800 8518 856
rect 8686 800 8702 856
rect 8870 800 8886 856
rect 9054 800 9070 856
rect 9238 800 9254 856
rect 9422 800 9438 856
rect 9606 800 9622 856
rect 9790 800 9806 856
rect 9974 800 9990 856
rect 10158 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10726 856
rect 10894 800 10910 856
rect 11078 800 11094 856
rect 11262 800 11278 856
rect 11446 800 11462 856
rect 11630 800 11646 856
rect 11814 800 11830 856
rect 11998 800 12014 856
rect 12182 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12566 856
rect 12734 800 12750 856
rect 12918 800 12934 856
rect 13102 800 13118 856
rect 13286 800 13302 856
rect 13470 800 13486 856
rect 13654 800 13670 856
rect 13838 800 13854 856
rect 14022 800 14038 856
rect 14206 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14590 856
rect 14758 800 14774 856
rect 14942 800 14958 856
rect 15126 800 15142 856
rect 15310 800 15326 856
rect 15494 800 15510 856
rect 15678 800 15694 856
rect 15862 800 15878 856
rect 16046 800 16062 856
rect 16230 800 16246 856
rect 16414 800 16430 856
rect 16598 800 16614 856
rect 16782 800 16798 856
rect 16966 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17350 856
rect 17518 800 17534 856
rect 17702 800 17718 856
rect 17886 800 17902 856
rect 18070 800 18086 856
rect 18254 800 18270 856
rect 18438 800 18454 856
rect 18622 800 18638 856
rect 18806 800 18822 856
rect 18990 800 19006 856
rect 19174 800 19190 856
rect 19358 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20110 856
rect 20278 800 20294 856
rect 20462 800 20478 856
rect 20646 800 20662 856
rect 20830 800 20846 856
rect 21014 800 21030 856
rect 21198 800 21214 856
rect 21382 800 21398 856
rect 21566 800 21582 856
rect 21750 800 21766 856
rect 21934 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22318 856
rect 22486 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22870 856
rect 23038 800 23054 856
rect 23222 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23790 856
rect 23958 800 23974 856
rect 24142 800 24158 856
rect 24326 800 24342 856
rect 24510 800 24526 856
rect 24694 800 24710 856
rect 24878 800 24894 856
rect 25062 800 25078 856
rect 25246 800 25262 856
rect 25430 800 25446 856
rect 25614 800 25630 856
rect 25798 800 25814 856
rect 25982 800 25998 856
rect 26166 800 26182 856
rect 26350 800 26366 856
rect 26534 800 26550 856
rect 26718 800 26734 856
rect 26902 800 26918 856
rect 27086 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27654 856
rect 27822 800 27838 856
rect 28006 800 28022 856
rect 28190 800 28206 856
rect 28374 800 28390 856
rect 28558 800 28574 856
rect 28742 800 28758 856
rect 28926 800 28942 856
rect 29110 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29494 856
rect 29662 800 29678 856
rect 29846 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30230 856
rect 30398 800 30414 856
rect 30582 800 30598 856
rect 30766 800 30782 856
rect 30950 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31334 856
rect 31502 800 31518 856
rect 31686 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32070 856
rect 32238 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32622 856
rect 32790 800 32806 856
rect 32974 800 32990 856
rect 33158 800 33174 856
rect 33342 800 33358 856
rect 33526 800 33542 856
rect 33710 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34094 856
rect 34262 800 34278 856
rect 34446 800 34462 856
rect 34630 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35198 856
rect 35366 800 35382 856
rect 35550 800 35566 856
rect 35734 800 35750 856
rect 35918 800 35934 856
rect 36102 800 36118 856
rect 36286 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36854 856
rect 37022 800 37038 856
rect 37206 800 37222 856
rect 37390 800 37406 856
rect 37574 800 37590 856
rect 37758 800 37774 856
rect 37942 800 37958 856
rect 38126 800 38142 856
rect 38310 800 38326 856
rect 38494 800 38510 856
rect 38678 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39062 856
rect 39230 800 39246 856
rect 39414 800 39430 856
rect 39598 800 39614 856
rect 39782 800 39798 856
rect 39966 800 39982 856
rect 40150 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40534 856
rect 40702 800 40718 856
rect 40886 800 40902 856
rect 41070 800 41086 856
rect 41254 800 41270 856
rect 41438 800 41454 856
rect 41622 800 41638 856
rect 41806 800 41822 856
rect 41990 800 42006 856
rect 42174 800 42190 856
rect 42358 800 42374 856
rect 42542 800 42558 856
rect 42726 800 42742 856
rect 42910 800 42926 856
rect 43094 800 43110 856
rect 43278 800 43294 856
rect 43462 800 43478 856
rect 43646 800 43662 856
rect 43830 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44398 856
rect 44566 800 44582 856
rect 44750 800 44766 856
rect 44934 800 44950 856
rect 45118 800 45134 856
rect 45302 800 45318 856
rect 45486 800 45502 856
rect 45670 800 45686 856
rect 45854 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46238 856
rect 46406 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46790 856
rect 46958 800 46974 856
rect 47142 800 47158 856
rect 47326 800 47342 856
rect 47510 800 47526 856
rect 47694 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48262 856
rect 48430 800 48446 856
rect 48614 800 48630 856
rect 48798 800 48814 856
rect 48982 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49550 856
rect 49718 800 49734 856
rect 49902 800 49918 856
rect 50086 800 50102 856
rect 50270 800 50286 856
rect 50454 800 50470 856
rect 50638 800 50654 856
rect 50822 800 50838 856
rect 51006 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51390 856
rect 51558 800 51574 856
rect 51742 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52126 856
rect 52294 800 52310 856
rect 52478 800 52494 856
rect 52662 800 52678 856
rect 52846 800 52862 856
rect 53030 800 53046 856
rect 53214 800 53230 856
rect 53398 800 53414 856
rect 53582 800 53598 856
rect 53766 800 53782 856
rect 53950 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54334 856
rect 54502 800 54518 856
rect 54686 800 54702 856
rect 54870 800 54886 856
rect 55054 800 55070 856
rect 55238 800 55254 856
rect 55422 800 55438 856
rect 55606 800 55622 856
rect 55790 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56174 856
rect 56342 800 56358 856
rect 56526 800 56542 856
rect 56710 800 56726 856
rect 56894 800 56910 856
rect 57078 800 57094 856
rect 57262 800 57278 856
rect 57446 800 57462 856
rect 57630 800 57646 856
rect 57814 800 57830 856
rect 57998 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58382 856
rect 58550 800 58566 856
rect 58734 800 58750 856
rect 58918 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59302 856
rect 59470 800 59486 856
rect 59654 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60038 856
rect 60206 800 60222 856
rect 60390 800 60406 856
rect 60574 800 60590 856
rect 60758 800 60774 856
rect 60942 800 60958 856
rect 61126 800 61142 856
rect 61310 800 61326 856
rect 61494 800 61510 856
rect 61678 800 61694 856
rect 61862 800 61878 856
rect 62046 800 62062 856
rect 62230 800 62246 856
rect 62414 800 62430 856
rect 62598 800 62614 856
rect 62782 800 62798 856
rect 62966 800 62982 856
rect 63150 800 63166 856
rect 63334 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63902 856
rect 64070 800 64086 856
rect 64254 800 64270 856
rect 64438 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64822 856
rect 64990 800 65006 856
rect 65174 800 65190 856
rect 65358 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66110 856
rect 66278 800 66294 856
rect 66462 800 66478 856
rect 66646 800 66662 856
rect 66830 800 66846 856
rect 67014 800 67030 856
rect 67198 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67582 856
rect 67750 800 67766 856
rect 67934 800 67950 856
rect 68118 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68686 856
rect 68854 800 68870 856
rect 69038 800 69054 856
rect 69222 800 69238 856
rect 69406 800 69422 856
rect 69590 800 69606 856
rect 69774 800 69790 856
rect 69958 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70342 856
rect 70510 800 70526 856
rect 70694 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71446 856
rect 71614 800 71630 856
rect 71798 800 71814 856
rect 71982 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72366 856
rect 72534 800 72550 856
rect 72718 800 72734 856
rect 72902 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73286 856
rect 73454 800 73470 856
rect 73638 800 73654 856
rect 73822 800 73838 856
rect 74006 800 74022 856
rect 74190 800 74206 856
rect 74374 800 74390 856
rect 74558 800 74574 856
rect 74742 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75310 856
rect 75478 800 75494 856
rect 75662 800 75678 856
rect 75846 800 75862 856
rect 76030 800 76046 856
rect 76214 800 76230 856
rect 76398 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76782 856
rect 76950 800 76966 856
rect 77134 800 77150 856
rect 77318 800 77334 856
rect 77502 800 77518 856
rect 77686 800 77702 856
rect 77870 800 77886 856
rect 78054 800 78070 856
rect 78238 800 78254 856
rect 78422 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78806 856
rect 78974 800 78990 856
rect 79158 800 79174 856
rect 79342 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79726 856
rect 79894 800 79910 856
rect 80078 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80646 856
rect 80814 800 80830 856
rect 80998 800 81014 856
rect 81182 800 81198 856
rect 81366 800 81382 856
rect 81550 800 81566 856
rect 81734 800 81750 856
rect 81918 800 81934 856
rect 82102 800 82118 856
rect 82286 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82854 856
rect 83022 800 83038 856
rect 83206 800 83222 856
rect 83390 800 83406 856
rect 83574 800 83590 856
rect 83758 800 83774 856
rect 83942 800 83958 856
rect 84126 800 84142 856
rect 84310 800 84326 856
rect 84494 800 84510 856
rect 84678 800 84694 856
rect 84862 800 84878 856
rect 85046 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85430 856
rect 85598 800 85614 856
rect 85782 800 85798 856
rect 85966 800 85982 856
rect 86150 800 86166 856
rect 86334 800 86350 856
rect 86518 800 86534 856
rect 86702 800 86718 856
rect 86886 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88006 856
rect 88174 800 88190 856
rect 88358 800 88374 856
rect 88542 800 88558 856
rect 88726 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89110 856
rect 89278 800 89294 856
rect 89462 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90214 856
rect 90382 800 90398 856
rect 90566 800 90582 856
<< obsm3 >>
rect 4208 2143 81328 90337
<< metal4 >>
rect 4208 2128 4528 90352
rect 19568 2128 19888 90352
rect 34928 2128 35248 90352
rect 50288 2128 50608 90352
rect 65648 2128 65968 90352
rect 81008 2128 81328 90352
<< labels >>
rlabel metal2 s 386 92026 442 92826 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24214 92026 24270 92826 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 26606 92026 26662 92826 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 28998 92026 29054 92826 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 31390 92026 31446 92826 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 33782 92026 33838 92826 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 36174 92026 36230 92826 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38566 92026 38622 92826 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40958 92026 41014 92826 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43350 92026 43406 92826 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45742 92026 45798 92826 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2686 92026 2742 92826 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 48042 92026 48098 92826 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50434 92026 50490 92826 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 52826 92026 52882 92826 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 55218 92026 55274 92826 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57610 92026 57666 92826 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 60002 92026 60058 92826 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 62394 92026 62450 92826 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 64786 92026 64842 92826 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 67178 92026 67234 92826 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 69570 92026 69626 92826 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5078 92026 5134 92826 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 71962 92026 72018 92826 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 74354 92026 74410 92826 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 76746 92026 76802 92826 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 79138 92026 79194 92826 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 81530 92026 81586 92826 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 83922 92026 83978 92826 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 86314 92026 86370 92826 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 88706 92026 88762 92826 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7470 92026 7526 92826 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 9862 92026 9918 92826 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12254 92026 12310 92826 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14646 92026 14702 92826 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17038 92026 17094 92826 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19430 92026 19486 92826 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 21822 92026 21878 92826 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1122 92026 1178 92826 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 25042 92026 25098 92826 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27434 92026 27490 92826 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29826 92026 29882 92826 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32126 92026 32182 92826 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34518 92026 34574 92826 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36910 92026 36966 92826 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39302 92026 39358 92826 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41694 92026 41750 92826 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 44086 92026 44142 92826 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46478 92026 46534 92826 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3514 92026 3570 92826 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48870 92026 48926 92826 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 51262 92026 51318 92826 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 53654 92026 53710 92826 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 56046 92026 56102 92826 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 58438 92026 58494 92826 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 60830 92026 60886 92826 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 63222 92026 63278 92826 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 65614 92026 65670 92826 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 68006 92026 68062 92826 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 70398 92026 70454 92826 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 5906 92026 5962 92826 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 72790 92026 72846 92826 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 75182 92026 75238 92826 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 77482 92026 77538 92826 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 79874 92026 79930 92826 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 82266 92026 82322 92826 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 84658 92026 84714 92826 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 87050 92026 87106 92826 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 89442 92026 89498 92826 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8298 92026 8354 92826 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10690 92026 10746 92826 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13082 92026 13138 92826 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15474 92026 15530 92826 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17866 92026 17922 92826 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20258 92026 20314 92826 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 22650 92026 22706 92826 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1950 92026 2006 92826 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 25778 92026 25834 92826 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28170 92026 28226 92826 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 30562 92026 30618 92826 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 32954 92026 33010 92826 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35346 92026 35402 92826 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37738 92026 37794 92826 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 40130 92026 40186 92826 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42522 92026 42578 92826 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44914 92026 44970 92826 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 47306 92026 47362 92826 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4342 92026 4398 92826 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 49698 92026 49754 92826 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 52090 92026 52146 92826 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 54482 92026 54538 92826 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 56874 92026 56930 92826 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 59266 92026 59322 92826 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 61566 92026 61622 92826 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 63958 92026 64014 92826 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 66350 92026 66406 92826 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 68742 92026 68798 92826 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 71134 92026 71190 92826 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6734 92026 6790 92826 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 73526 92026 73582 92826 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 75918 92026 75974 92826 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 78310 92026 78366 92826 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 80702 92026 80758 92826 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 83094 92026 83150 92826 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 85486 92026 85542 92826 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 87878 92026 87934 92826 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 90270 92026 90326 92826 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9126 92026 9182 92826 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11518 92026 11574 92826 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 13910 92026 13966 92826 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16210 92026 16266 92826 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18602 92026 18658 92826 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 20994 92026 21050 92826 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23386 92026 23442 92826 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 90352 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 90352 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 90352 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 90352 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 90352 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 90352 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 90682 92826
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 13448332
string GDS_START 245544
<< end >>

